**.subckt untitled-1
x1 GND p1 lc
V1 p1 GND 3
**** begin user architecture code

.ac lin 10k 1G 5G
.end
.control
destroy all
run
plot i(v1)
plot v(v1)
plot v(v1)/i(v1)
.endc

**** end user architecture code
**.ends

* expanding   symbol:  lc.sym # of pins=2
* sym_path: /home/hugodg/projects_sky130/microelectronic/LC/xschem/lc.sym
* sch_path: /home/hugodg/projects_sky130/microelectronic/LC/xschem/lc.sch
.subckt lc  p2 p1
*.iopin p1
*.iopin p2
L1 p1 p2 5.092n m=3
C1 p1 p2 828.74f m=1
.ends

.GLOBAL GND
.end
