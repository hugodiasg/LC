magic
tech sky130A
timestamp 1639090007
<< metal4 >>
rect 4400 12979 5200 19300
rect 4400 12221 4420 12979
rect 5178 12221 5200 12979
rect 4400 12200 5200 12221
<< via4 >>
rect 4420 12221 5178 12979
<< metal5 >>
rect 0 17700 18500 18500
rect 0 16600 17400 17400
rect 0 800 800 16600
rect 1100 15500 16300 16300
rect 1100 1900 1900 15500
rect 2200 14400 15200 15200
rect 2200 3000 3000 14400
rect 3300 13300 14100 14100
rect 3300 4100 4100 13300
rect 4400 12979 5200 13000
rect 4400 12221 4420 12979
rect 5178 12221 5200 12979
rect 4400 5200 5200 12221
rect 13300 5200 14100 13300
rect 4400 4400 14100 5200
rect 14400 4100 15200 14400
rect 3300 3300 15200 4100
rect 15500 3000 16300 15500
rect 2200 2200 16300 3000
rect 16600 1900 17400 16600
rect 1100 1100 17400 1900
rect 17700 800 18500 17700
rect 0 0 18500 800
<< end >>
