magic
tech sky130A
magscale 1 2
timestamp 1638043154
<< metal4 >>
rect -9022 47378 -3022 53378
rect -6938 45008 -5338 47378
rect -15446 43414 10408 45008
rect -15446 39516 -13846 43414
rect -2810 43408 10408 43414
rect -35872 36730 -13846 39516
rect 8808 38992 10408 43408
rect 8808 38486 10412 38992
rect -35872 17516 -13872 36730
<< metal5 >>
rect -35872 38398 -13872 39516
rect -35872 36798 3706 38398
rect -35872 17516 -13872 36798
rect -7018 33760 -5418 36798
rect -9188 27760 -3188 33760
use 1  1_0
timestamp 1638042750
transform 1 0 98 0 1 -23
box 0 0 38400 40000
<< labels >>
flabel metal5 -6240 30430 -6240 30430 0 FreeSans 32000 0 0 0 P1
flabel metal4 -5956 50414 -5956 50414 0 FreeSans 32000 0 0 0 P2
<< end >>
