magic
tech sky130A
timestamp 1638042750
<< metal4 >>
rect 4400 13679 5200 20000
rect 4400 12921 4420 13679
rect 5178 12921 5200 13679
rect 4400 12900 5200 12921
<< via4 >>
rect 4420 12921 5178 13679
<< metal5 >>
rect 0 18400 19200 19200
rect 0 17300 18100 18100
rect 0 800 800 17300
rect 1100 16200 17000 17000
rect 1100 1900 1900 16200
rect 2200 15100 15900 15900
rect 2200 3000 3000 15100
rect 3300 14000 14800 14800
rect 3300 4100 4100 14000
rect 4400 13679 5200 13700
rect 4400 12921 4420 13679
rect 5178 12921 5200 13679
rect 4400 5200 5200 12921
rect 14000 5200 14800 14000
rect 4400 4400 14800 5200
rect 15100 4100 15900 15100
rect 3300 3300 15900 4100
rect 16200 3000 17000 16200
rect 2200 2200 17000 3000
rect 17300 1900 18100 17300
rect 1100 1100 18100 1900
rect 18400 800 19200 18400
rect 0 0 19200 800
<< end >>
