magic
tech sky130A
magscale 1 2
timestamp 1639092644
<< metal3 >>
rect 12400 23800 14300 24000
rect 12400 22600 12700 23800
rect 13900 22600 14300 23800
rect 12400 8100 14300 22600
rect 12400 6400 17500 8100
rect 12400 4400 14300 6400
rect 12400 4100 13200 4400
rect 15800 100 17500 6400
rect 15800 -13000 17600 100
<< via3 >>
rect 12700 22600 13900 23800
<< metal4 >>
rect 9200 24700 28900 26100
rect 10600 4100 11700 24700
rect 27900 24500 28900 24700
rect 12699 23800 13901 23801
rect 12699 22600 12700 23800
rect 13900 22600 13901 23800
rect 12699 22599 13901 22600
<< via4 >>
rect 12700 22600 13900 23800
<< metal5 >>
rect 12400 23800 40600 24000
rect 12400 22600 12700 23800
rect 13900 22600 40600 23800
rect 12400 22400 40600 22600
use sky130_fd_pr__cap_mim_m3_1_NUZ66F  XC0
timestamp 1639088392
transform 1 0 12367 0 1 2517
box -2167 -2117 2166 2117
use l0  l0_0
timestamp 1639090007
transform 1 0 18523 0 1 -12908
box 0 0 37000 38600
<< labels >>
flabel metal4 9500 25000 10300 25900 0 FreeSans 1600 0 0 0 p1
port 1 nsew
flabel metal3 16300 -12700 17300 -11700 0 FreeSans 1600 0 0 0 p2
port 2 nsew
<< end >>
